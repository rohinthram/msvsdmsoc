* SPICE3 file created from inverter.ext - technology: sky130A

.lib ~/Downloads/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option scale=10000u

X0 out in vdd w_n192_142# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=98 l=30
X1 out in vss SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=98 l=30

v1 vdd gnd dc 1
v2 vss gnd dc -1

v3 in gnd PULSE(-1 1 0 0 0 1u 2u)

.tran 0.1u 10u

.control
run
plot v(out)
plot v(in)
.endc

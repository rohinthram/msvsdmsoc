* SPICE3 file created from inverter.ext - technology: sky130A

.option scale=10000u

X0 out in vdd w_n192_142# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=98 l=30
X1 out in vss SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=98 l=30
